


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity RECV_RPM is
 Port ( 
    RPM
 );
end RECV_RPM;

architecture Behavioral of RECV_RPM is

begin


end Behavioral;
